interface IfMEM();

    wire        dqs_p;
    wire        dqs_n;
    wire        dq;

endinterface